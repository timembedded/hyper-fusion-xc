-- 
-- VoiceRom.vhd 
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.VM2413.ALL;

entity VoiceRom is 
  port (  
    clk    : in std_logic;
    addr : in VOICE_ID_TYPE;
    data  : out VOICE_TYPE
  );
end VoiceRom;

architecture RTL of VoiceRom is

  type VOICE_ARRAY_TYPE is array (VOICE_ID_TYPE'range) of VOICE_VECTOR_TYPE;
  constant voices : VOICE_ARRAY_TYPE := (
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "0" & "0" & "0000" & "00" & "000000" & "0" & "000" & "0000" & "0000" & "0000" & "0000", -- @0(M)
  "0" & "0" & "0" & "0" & "0000" & "00" & "000000" & "0" & "000" & "0000" & "0000" & "0000" & "0000", -- @0(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "1" & "1" & "0" & "0001" & "00" & "011110" & "0" & "111" & "1111" & "0000" & "0000" & "0000", -- @1(M)
  "0" & "1" & "1" & "0" & "0001" & "00" & "000000" & "1" & "000" & "0111" & "1111" & "0001" & "0111", -- @1(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "0" & "1" & "0011" & "00" & "010111" & "1" & "110" & "1111" & "1111" & "0010" & "0011", -- @2(M)
  "0" & "1" & "0" & "0" & "0001" & "00" & "000000" & "0" & "000" & "1111" & "1111" & "0001" & "0011", -- @2(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0011" & "10" & "011010" & "0" & "100" & "1010" & "0011" & "1111" & "0000", -- @3(M)
  "0" & "0" & "0" & "0" & "0001" & "00" & "000000" & "0" & "000" & "1111" & "0100" & "0010" & "0011", -- @3(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "0" & "1" & "0001" & "00" & "001110" & "0" & "111" & "1111" & "1010" & "0111" & "0000", -- @4(M)
  "0" & "1" & "1" & "0" & "0001" & "00" & "000000" & "0" & "000" & "0110" & "0100" & "0001" & "0111", -- @4(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0010" & "00" & "011110" & "0" & "110" & "1111" & "0000" & "0000" & "0000", -- @5(M)
  "0" & "0" & "1" & "0" & "0001" & "00" & "000000" & "0" & "000" & "0111" & "0110" & "0010" & "1000", -- @5(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0001" & "00" & "010110" & "0" & "101" & "1111" & "0000" & "0000" & "0000", -- @6(M)
  "0" & "0" & "1" & "0" & "0010" & "00" & "000000" & "0" & "000" & "0111" & "0001" & "0001" & "1000", -- @6(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0001" & "00" & "011101" & "0" & "111" & "1000" & "0010" & "0001" & "0000", -- @7(M)
  "0" & "1" & "1" & "0" & "0001" & "00" & "000000" & "0" & "000" & "1000" & "0000" & "0000" & "0111", -- @7(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0011" & "00" & "101101" & "0" & "110" & "1001" & "0000" & "0000" & "0000", -- @8(M)
  "0" & "0" & "1" & "0" & "0001" & "00" & "000000" & "1" & "000" & "1001" & "0000" & "0000" & "0111", -- @8(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0001" & "00" & "011011" & "0" & "110" & "0110" & "0100" & "0001" & "0000", -- @9(M)
  "0" & "0" & "1" & "0" & "0001" & "00" & "000000" & "0" & "000" & "0110" & "0101" & "0001" & "0111", -- @9(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0001" & "00" & "001011" & "1" & "010" & "1000" & "0101" & "0111" & "0000", -- @10(M)
  "0" & "0" & "1" & "0" & "0001" & "00" & "000000" & "1" & "000" & "1010" & "0000" & "0000" & "0111", -- @10(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0011" & "10" & "000011" & "0" & "000" & "1111" & "1111" & "0001" & "0000", -- @11(M)
  "0" & "0" & "0" & "0" & "0001" & "00" & "000000" & "1" & "000" & "1011" & "0000" & "0000" & "0100", -- @11(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "1" & "0" & "0" & "1" & "0111" & "00" & "100000" & "0" & "111" & "1111" & "1111" & "0010" & "0010", -- @12(M)
  "1" & "1" & "0" & "0" & "0001" & "00" & "000000" & "0" & "000" & "1111" & "1111" & "0001" & "0010", -- @12(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "1" & "1" & "0" & "0001" & "00" & "001100" & "0" & "101" & "1101" & "0010" & "0100" & "0000", -- @13(M)
  "0" & "0" & "0" & "0" & "0000" & "00" & "000000" & "0" & "000" & "1111" & "0110" & "0100" & "0011", -- @13(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "0" & "0" & "0001" & "01" & "010110" & "0" & "011" & "1111" & "0100" & "0000" & "0011", -- @14(M)
  "0" & "0" & "0" & "0" & "0001" & "00" & "000000" & "0" & "000" & "1111" & "0000" & "0000" & "0010", -- @14(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0001" & "10" & "001001" & "0" & "011" & "1111" & "0001" & "1111" & "0000", -- @15(M)
  "0" & "1" & "0" & "0" & "0001" & "00" & "000000" & "0" & "000" & "1111" & "0100" & "0010" & "0011", -- @15(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "0" & "0" & "0111" & "00" & "010110" & "0" & "000" & "1101" & "1111" & "1111" & "1111", -- BD(M)
  "0" & "0" & "1" & "0" & "0001" & "00" & "000000" & "0" & "000" & "1111" & "1000" & "1111" & "1000", -- BD(C)
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "1" & "0001" & "00" & "000000" & "0" & "000" & "1111" & "0111" & "1111" & "0111", -- HH
  "0" & "0" & "1" & "1" & "0010" & "00" & "000000" & "0" & "000" & "1111" & "0111" & "1111" & "0111", -- SD
-- AM    PM    EG    KR     ML      KL       TL       WF    FB       AR       DR       SL       RR
  "0" & "0" & "1" & "0" & "0101" & "00" & "000000" & "0" & "000" & "1111" & "1000" & "1111" & "1000", -- TOM
  "0" & "0" & "0" & "0" & "0001" & "00" & "000000" & "0" & "000" & "1101" & "1100" & "0101" & "0101"  -- CYM
);

begin

  process (clk) 

  begin
  
    if clk'event and clk = '1' then
	  data <= CONV_VOICE(voices(addr));
    end if;
    
  end process;

end RTL;